`include "../src/RTL/define.v"
`define   CYCLE   8
`define   TOTAL_CYCLE 50000
`timescale 1ns/100ps


module tb;

reg                       sys_clk;
reg                       sys_rst;

reg   [`WIDTH-1:0]        CPU0_instruction;
reg   [`WIDTH-1:0]        CPU0_write_data_i;
                     
wire                      CPU0_data_en_o;
wire  [`WIDTH-1:0]        CPU0_read_data_o;
                     
reg   [`WIDTH-1:0]        CPU1_instruction;
reg   [`WIDTH-1:0]        CPU1_write_data_i;
                     
wire                      CPU1_data_en_o;
wire  [`WIDTH-1:0]        CPU1_read_data_o;

reg   [4:0]               error_num;
reg   [4:0]               counter;


top top_SoC (
    .sys_clk            (sys_clk),
    .sys_rst            (sys_rst),

    .CPU0_instruction   (CPU0_instruction),
    .CPU0_write_data_i  (CPU0_write_data_i), 

    .CPU0_data_en_o     (CPU0_data_en_o),
    .CPU0_read_data_o   (CPU0_read_data_o),
 
    .CPU1_instruction   (CPU1_instruction),
    .CPU1_write_data_i  (CPU1_write_data_i),
    
    .CPU1_data_en_o     (CPU1_data_en_o),
    .CPU1_read_data_o   (CPU1_read_data_o) 
);

always begin
    #(`CYCLE/2) sys_clk = ~sys_clk;
end


initial begin
    sys_clk   = 0;
    sys_rst   = 1;
    

    #(`CYCLE);
    sys_rst   = 0;
    #(`CYCLE/2)
    error_num = 0;
    counter   = 0;
    
    
    
    /**********************************************************************
                         Local CPU READ WRITE TEST
    **********************************************************************/
    
    
    
    /**********************************************************************
        1. 
            CPU0 / write / miss / sw x5, 0(x0)
            id   : 0
            tag  : 0
            data : 1010_1010
            state: I -> M
    **********************************************************************/
    CPU0_instruction = 32'h00502023;
    CPU0_write_data_i = 32'h1010_1010;
    counter = counter + 1;
    #(`CYCLE); 
    CPU0_instruction = 32'h0;

    wait(CPU0_data_en_o);
    #(`CYCLE*2);
    $display("1.  CPU0 write, id = 0, tag = 0, write data = 1010_1010 / M");
    
    
    /**********************************************************************
        2. 
            CPU0 / write / hit / sw x5, 0(x0)
            id   : 0
            tag  : 0
            data : 2020_2020
            state: M -> M
    **********************************************************************/    
    CPU0_instruction = 32'h00502023;
    CPU0_write_data_i = 32'h2020_2020;
    counter = counter + 1;
    #(`CYCLE); 
    CPU0_instruction = 32'h0;

    wait(CPU0_data_en_o);
    #(`CYCLE*2);
    $display("2.  CPU0 write, id = 0, tag = 0, write data = 2020_2020 / M");

    /**********************************************************************
        3. 
            CPU0 / read / hit / lw x5, 0(x0)
            id   : 0
            tag  : 0
            data : 2020_2020
            state: M -> M
    **********************************************************************/      
    CPU0_instruction = 32'h00002283;
    counter = counter + 1;
    #(`CYCLE); 
    CPU0_instruction = 32'h0;

    wait(CPU0_data_en_o);
    #(`CYCLE*2);
    if (CPU0_read_data_o != 32'h2020_2020) begin
        error_num = error_num + 1;
    end
    $display("3.  CPU0 read,  id = 0, tag = 0, read  data = %h (expect: 2020_2020)/ M", CPU0_read_data_o);    
    

    /**********************************************************************
        4. 
            CPU0 / read / miss / lw x5, 256(x0)
            id   : 0
            tag  : 1
            data : 1
            state: I -> E
    **********************************************************************/       
    CPU0_instruction = 32'h10002283;
    counter = counter + 1;
    #(`CYCLE); 
    CPU0_instruction = 32'h0;

    wait(CPU0_data_en_o);
    #(`CYCLE*2);
    if (CPU0_read_data_o != 32'h1) begin
        error_num = error_num + 1;
    end
    $display("4.  CPU0 read,  id = 0, tag = 1, read  data = %h (expect: 1)/ E", CPU0_read_data_o);  
    

    /**********************************************************************
        5. 
            CPU0 / read / hit / lw x5, 256(x0)
            id   : 0
            tag  : 1
            data : 1
            state: E -> E
    **********************************************************************/       
    CPU0_instruction = 32'h10002283; 
    counter = counter + 1;
    #(`CYCLE); 
    CPU0_instruction = 32'h0;

    wait(CPU0_data_en_o);
    #(`CYCLE*2);
    if (CPU0_read_data_o != 32'h1) begin
        error_num = error_num + 1;
    end
    $display("5.  CPU0 read,  id = 0, tag = 1, read  data = %h (expect: 1)/ E", CPU0_read_data_o);  
    
    
    /**********************************************************************
        6. 
            CPU0 / write / hit / sw x5, 256(x0)
            id   : 0
            tag  : 1
            data : 3030_3030
            state: E -> M
    **********************************************************************/    
    CPU0_instruction = 32'h10502023; // sw x5, 32(x0)
    CPU0_write_data_i = 32'h3030_3030;
    counter = counter + 1;
    #(`CYCLE); 
    CPU0_instruction = 32'h0;

    wait(CPU0_data_en_o);
    #(`CYCLE*2);
    $display("6.  CPU0 write, id = 0, tag = 1, write data = 3030_3030 / M"); 


    /**********************************************************************
        7. 
            CPU0 / read / miss / lw x5, 512(x0)
            id   : 0
            tag  : 2
            data : 1
            state: I -> E
    **********************************************************************/     
    CPU0_instruction = 32'h20002283; 
    counter = counter + 1;
    #(`CYCLE); 
    CPU0_instruction = 32'h0;

    wait(CPU0_data_en_o);
    #(`CYCLE*2);
    if (CPU0_read_data_o != 32'h1) begin
        error_num = error_num + 1;
    end
    $display("7.  CPU0 read,  id = 0, tag = 2, read  data = %h (expect: 1)/ E", CPU0_read_data_o);

    /**********************************************************************
        8. 
            CPU0 / read / miss / lw x5, 768(x0)
            id   : 0
            tag  : 3
            data : 1
            state: I -> E
    **********************************************************************/      
    CPU0_instruction = 32'h30002283;
    counter = counter + 1;
    #(`CYCLE); 
    CPU0_instruction = 32'h0;

    wait(CPU0_data_en_o);
    #(`CYCLE*2);
    if (CPU0_read_data_o != 32'h1) begin
        error_num = error_num + 1;
    end
    $display("8.  CPU0 read,  id = 0, tag = 3, read  data = %h (expect: 1)/ E", CPU0_read_data_o);    






    /**********************************************************************
                              FORWARD TEST
    **********************************************************************/

    /**********************************************************************
        9. 
            CPU1 / read / miss / lw x5, 0(x0)
            id   : 0
            tag  : 0
            data : 2020_2020
            state: I -> S, state': M -> S
    **********************************************************************/      
    CPU1_instruction = 32'h00002283;
    counter = counter + 1;
    #(`CYCLE); 
    CPU1_instruction = 32'h0;

    wait(CPU1_data_en_o);
    #(`CYCLE*2);
    if (CPU1_read_data_o != 32'h2020_2020) begin
        error_num = error_num + 1;
    end
    $display("9.  CPU1 read,  id = 0, tag = 0, read  data = %h (expect: 2020_2020)/ S", CPU1_read_data_o); 

    /**********************************************************************
        10. 
            CPU1 / read / hit / lw x5, 0(x0)
            id   : 0
            tag  : 0
            data : 2020_2020
            state: S -> S, state': S -> S
    **********************************************************************/      
    CPU1_instruction = 32'h00002283;
    counter = counter + 1;
    #(`CYCLE); 
    CPU1_instruction = 32'h0;

    wait(CPU1_data_en_o);
    #(`CYCLE*2);
    if (CPU1_read_data_o != 32'h2020_2020) begin
        error_num = error_num + 1;
    end
    $display("10. CPU1 read,  id = 0, tag = 0, read  data = %h (expect: 2020_2020)/ S", CPU1_read_data_o);      
    
    /**********************************************************************
        11. 
            CPU1 / write / hit / sw x5, 0(x0)
            id   : 0
            tag  : 0
            data : 4040_4040
            state: S -> M, state': S -> I
    **********************************************************************/
    CPU1_instruction = 32'h00502023;
    CPU1_write_data_i = 32'h4040_4040;
    counter = counter + 1;
    #(`CYCLE); 
    CPU1_instruction = 32'h0;

    wait(CPU1_data_en_o);
    #(`CYCLE*2);
    $display("11. CPU1 write, id = 0, tag = 0, write data = 4040_4040 / M");    
    
    /**********************************************************************
        12. 
            CPU1 / write / miss / sw x5, 256(x0)
            id   : 0
            tag  : 1
            data : 5050_5050
            state: I -> M, state': M -> I
    **********************************************************************/
    CPU1_instruction = 32'h10502023;
    CPU1_write_data_i = 32'h5050_5050;
    counter = counter + 1;
    #(`CYCLE); 
    CPU1_instruction = 32'h0;

    wait(CPU1_data_en_o);
    #(`CYCLE*2);
    $display("11. CPU1 write, id = 0, tag = 1, write data = 5050_5050 / M");  

    /**********************************************************************
        13. 
            CPU1 / read / miss / lw x5, 512(x0)
            id   : 0
            tag  : 2
            data : 1
            state: I -> S, state': E -> S
    **********************************************************************/      
    CPU1_instruction = 32'h20002283;
    counter = counter + 1;
    #(`CYCLE); 
    CPU1_instruction = 32'h0;

    wait(CPU1_data_en_o);
    #(`CYCLE*2);
    if (CPU1_read_data_o != 32'h1) begin
        error_num = error_num + 1;
    end
    $display("13. CPU1 read,  id = 0, tag = 2, read  data = %h (expect: 1)/ S", CPU1_read_data_o);        
    
    /**********************************************************************
        14. 
            CPU1 / write / miss / sw x5, 768(x0)
            id   : 0
            tag  : 3
            data : 6060_6060
            state: I -> M, state': E -> I
    **********************************************************************/
    CPU1_instruction = 32'h30502023;
    CPU1_write_data_i = 32'h6060_6060;
    counter = counter + 1;
    #(`CYCLE); 
    CPU1_instruction = 32'h0;

    wait(CPU1_data_en_o);
    #(`CYCLE*2);
    $display("14. CPU1 write, id = 0, tag = 3, write data = 6060_6060 / M"); 
    
    /**********************************************************************
        15. 
            CPU0 / read / miss / lw x5, 768(x0)
            id   : 0
            tag  : 3
            data : 6060_6060
            state: I -> S, state': M -> S
    **********************************************************************/      
    CPU0_instruction = 32'h30002283;
    counter = counter + 1;
    #(`CYCLE); 
    CPU0_instruction = 32'h0;

    wait(CPU0_data_en_o);
    #(`CYCLE*2);
    if (CPU0_read_data_o != 32'h6060_6060) begin
        error_num = error_num + 1;
    end
    $display("15. CPU0 read,  id = 0, tag = 3, read  data = %h (expect: 6060_6060)/ S", CPU0_read_data_o);   
    
    /**********************************************************************
        16. 
            CPU1 / read / hit / lw x5, 768(x0)
            id   : 0
            tag  : 3
            data : 6060_6060
            state: S -> S, state': S -> S
    **********************************************************************/      
    CPU1_instruction = 32'h30002283;
    counter = counter + 1;
    #(`CYCLE); 
    CPU1_instruction = 32'h0;

    wait(CPU1_data_en_o);
    #(`CYCLE*2);
    if (CPU1_read_data_o != 32'h6060_6060) begin
        error_num = error_num + 1;
    end
    $display("16. CPU1 read,  id = 0, tag = 3, read  data = %h (expect: 6060_6060)/ S", CPU1_read_data_o);  

    /**********************************************************************
        17. 
            CPU1 / write / hit / sw x5, 512(x0)
            id   : 0
            tag  : 2
            data : 7070_7070
            state: S -> M, state': S -> I
    **********************************************************************/
    CPU1_instruction = 32'h20502023;
    CPU1_write_data_i = 32'h7070_7070;
    counter = counter + 1;
    #(`CYCLE); 
    CPU1_instruction = 32'h0;

    wait(CPU1_data_en_o);
    #(`CYCLE*2);
    $display("17. CPU1 write, id = 0, tag = 2, write data = 7070_7070 / M");  
    


    /**********************************************************************
                            LRU Replacement
    **********************************************************************/
   
    /**********************************************************************
        18. 
            CPU0 / write / miss / sw x5, 832(x0)
            id   : 1
            tag  : 2
            data : 8080_8080
            state: I -> M
    **********************************************************************/
    CPU0_instruction = 32'h24002283;
    CPU0_write_data_i = 32'h8080_8080;
    counter = counter + 1;
    #(`CYCLE); 
    CPU0_instruction = 32'h0;

    wait(CPU0_data_en_o);
    #(`CYCLE*2);
    $display("18. CPU0 write, id = 1, tag = 4, write data = 8080_8080 / M");  

    /**********************************************************************
        19. 
            CPU0 / write / miss / sw x5, 1088(x0)
            id   : 1
            tag  : 4
            data : 9090_9090
            state: I -> M
    **********************************************************************/
    CPU0_instruction = 32'h44502023;
    CPU0_write_data_i = 32'h9090_9090;
    counter = counter + 1;
    #(`CYCLE); 
    CPU0_instruction = 32'h0;

    wait(CPU0_data_en_o);
    #(`CYCLE*2);
    $display("19. CPU0 write, id = 1, tag = 4, write data = 9090_9090 / M");        
    
    /**********************************************************************
        20. 
            CPU0 / write / miss / sw x5, 1344(x0)
            id   : 1
            tag  : 5
            data : A0A0_A0A0
            state: I -> M
    **********************************************************************/
    CPU0_instruction = 32'h54502023;
    CPU0_write_data_i = 32'hA0A0_A0A0;
    counter = counter + 1;
    #(`CYCLE); 
    CPU0_instruction = 32'h0;

    wait(CPU0_data_en_o);
    #(`CYCLE*2);
    $display("20. CPU0 write, id = 1, tag = 6, write data = A0A0_A0A0 / M");      
    
    /**********************************************************************
        21. 
            CPU0 / write / miss / sw x5, 1600(x0)
            id   : 1
            tag  : 6
            data : B0B0_B0B0
            state: I -> M
    **********************************************************************/
    CPU0_instruction = 32'h64502023;
    CPU0_write_data_i = 32'hB0B0_B0B0;
    counter = counter + 1;
    #(`CYCLE); 
    CPU0_instruction = 32'h0;

    wait(CPU0_data_en_o);
    #(`CYCLE*2);
    $display("21. CPU0 write, id = 1, tag = 7, write data = B0B0_B0B0 / M"); 

    /**********************************************************************
        22. 
            CPU0 / write / miss / sw x5, 1856(x0)
            id   : 1
            tag  : 7
            data : C0C0_C0C0
            state: I -> M
    **********************************************************************/
    CPU0_instruction = 32'h74502023;
    CPU0_write_data_i = 32'hC0C0_C0C0;
    counter = counter + 1;
    #(`CYCLE); 
    CPU0_instruction = 32'h0;

    wait(CPU0_data_en_o);
    #(`CYCLE*2);
    $display("22. CPU0 write, id = 1, tag = 8, write data = C0C0_C0C0 / M");      

    /**********************************************************************
        23. 
            CPU0 / read / hit / lw x5, 1856(x0)
            id   : 1
            tag  : 7
            data : 1
            state: M -> M
    **********************************************************************/     
    CPU0_instruction = 32'h74002283; 
    counter = counter + 1;
    #(`CYCLE); 
    CPU0_instruction = 32'h0;

    wait(CPU0_data_en_o);
    #(`CYCLE*2);
    if (CPU0_read_data_o != 32'hC0C0_C0C0) begin
        error_num = error_num + 1;
    end
    $display("23. CPU0 read,  id = 1, tag = 8, read  data = %h (expect: C0C0_C0C0)/ M", CPU0_read_data_o); 

    
    if (error_num == 0) begin
        $display("");   
        $display("        ,@@@@@@@@@@,,@@@@@@@&  .#&@@@&&.,@@@@@@@@@@,      &@@@@@@&*   ,@@@&     .#&@@@&&.  *&@@@@&(  ,@@@@@@@&  &@@@@@,     ,@@,");
        $display("            ,@@,    ,@@,      ,@@/   ./.    ,@@,          &@&   ,&@# .&@&@@(   .@@/   ./. #@&.  .,/  ,@@,       &@&  *&@&.  ,@@,");
        $display("            ,@@,    ,@@&&&&&. .&@@/,        ,@@,          &@&   ,&@# &@& /@@,  .&@@/,     (@@&&(*.   ,@@&&&&&.  &@&    &@#  ,@@,");
        $display("            ,@@,    ,@@&&&&&. .&@@/,        ,@@,          &@&   ,&@# &@& /@@,  .&@@/,     (@@&&(*.   ,@@&&&&&.  &@&    &@#  ,@@,");
        $display("            ,@@,    ,@@/,,,,    ./#&@@@(    ,@@,          &@@@@@@&* /@@,  #@&.   ./#&@@@(   *(&&@@&. ,@@/,,,,   &@&    &@#  .&&.");
        $display("            ,@@,    ,@@,      ./,   .&@#    ,@@,          &@&      ,@@@@@@@@@& ./.   .&@# /*.   /@@. ,@@,       &@&  *&@&.   ,, ");
        $display("            ,@@,    ,@@@@@@@& .#&@@@@&/     ,@@,          &@&     .&@#     ,@@/.#&@@@@&/   /&&@@@@.  ,@@@@@@@&  &@@@@@.     ,@@,");
        $display(",*************,,*/(((((//,,*(#&&&&&&&&&&&&&&&#(*,,,****************************************************,*/(((((((((/((((////****/((##&&&&&&");
        $display(",*************,,//((((((//,,*(&&&&&&&&&&&&&&&&&##/*****************************************************,,*/(///(//////****//((##&&&&&&&&&&&");
        $display(",************,,*/(((((((//***/#&&&&&&&&&&&&&&&&&&&#(/***************************************************,*//////////*//((#&&&&&&&&&&&&&&&&&");
        $display(",***********,,*////////////***/##&&&&&&&&&&&&&&&&&&&##(*,***********************************************,,*////////(###&&&&&&&&&&&&&&&&&&&&");
        $display(",**********,,,*/*******//////**/(#&&&&&&&&&&&&&&&&&&&&&#(/**********************************************,,,***/(##&&&&&&&&&&&&&&&&&&&&&&&&&");
        $display(",*********,,,,*************///***/(#&&&&&&&&&&&&&&&&&&&&&&#(/***********************************,****,****/((#&&&&&&&&&&&&&&&&&&&&&&&&&&&&#");
        $display(",*********,,,***************//****/(##&&&&&&&&&&&&&&&&&&&&&&##//**************//////////////////////((#####&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&#(");
        $display(",********,,,,***********************/(#&&&&&&&&&&&&&&&&&&&&&&&##################&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&##(/");
        $display(",*******,..,***********************,,*/##&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&###((//");
        $display(",*******,.,,***********************,,,,*(#&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&##(//**//");
        $display(",******,.,,,************************,,,,*/(#&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&#(//*******");
        $display(",*****,,,,,********,***,,,,,,,,,,,,*,,,,,,*/(######&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&##(/**********");
        $display(",*****,..,*******,,,,,,,,,,,,,,,,,,,,,,*,,,,*///((#&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&###(/************");
        $display(",*****,,,*******,,,,,*,,,,,,,,,,,,,,,,,****,,,*/(#&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&#######(//**************");
        $display(",****,.,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,**,,,/(&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&#((//******************");
        $display(",***,..,,,,,,,,,,,,,,,,,,,,,,,,,,,,,..,,,,,,,*(#&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&#(/*******************");
        $display(",**,,.,,,,,,,,,,,,,,,,,,,,,,,,,,.......,,,,,,/#&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&#####&&&&&&&&&&&&&&&&#(/******************");
        $display(",**,..,,,,,,,,,,,,,,,,,,,,,,,,,......,,,*,,,*(#&&&&&&&&##(((/(##&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&##(((/*/((#&&&&&&&&&&&&&&#(/*****************");
        $display(",*,..,,,,,,,,,,,,,,,,,,,,,,,,,,,.....,,**,,*/#&&&&&&&##((((*,**/#&&&&&&&&&&&&&&&&&&&&&&&&&&&&##((##/,,,*(#&&&&&&&&&&&&&&#(*****************");
        $display(".*,.,,,**,,,,,,,,,,,,,,,,,,,,,,,,,,*****,,,/(&&&&&&&&#(//(#/,..*/#&&&&&&&&&&&&&&&&&&&&&&&&&&&#(//(#/,..,/(#&&&&&&&&&&&&&&#/*****///////////");
        $display(".,..,,,,,,,,,,,,,,,,,,,,,,,,,,*,,*******,,,(#&&&&&&&&#(*,,,....,/#&&&&&&&&&&&&&&&&&&&&&&&&&&&#(*,,,....,/(#&&&&&&&&&&&&&&#(*,**////////////");
        $display(".,..,,,,,,,,,...........,,,,,,*,********,,*(#&&&&&&&&&#(/*,,...,/#&&&&&&&&&&&&&&&&&&&&&&&&&&&&#(/*,,..,*/##&&&&&&&&&&&&&&&#(***////////////");
        $display(" ..,,,,,,.................,,,**********,,*(#&&&&&&&&&&&&&&&&&&#&&&&&&&&#((///((#&&&&&&&&&&&&&&&&&&&&&#&&&&&&&&&&&&&&&&&&&&&#/**////////////");
        $display(".,,,,,,,,.................,,***********,,/(####&&&&&&&&&&&&&&&&&&&&&&&&#(/*,,,*(#&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&#(/*////////////");
        $display(".,***,,,,,,..............,,,**********,..,***//((##&&&&&&&&&&&&&&&&&&&&&&&##((##&&&&&&&&&&&&&&&&&&&&&&&&&##(((((((((###&&&&&#/**///////////");
        $display(".*****,,,,,,,,,,,,,,,,,,,*************,..,*******/(#&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&##///*//////((#&&&&&#(**///////////");
        $display(".****************/******/***////*****,.,*///////**/#&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&#(////////////(#&&&&&#/**//////////");
        $display(".***********************/////*******,..,*//////////(#&&&&&&&&&&&&&&&&&&&&##########&&&&&&&&&&&&&&&&&&&&#(///////////*/(#&&&&&#(***/////////");
        $display(".************************///********,..,*//////////#&&&&&&&&&&&&&&&&&&#(//*****///(((##&&&&&&&&&&&&&&&&#(///////////**/##&&&&##/***////////");
        $display(".***********************************,.,,***///////(#&&&&&&&&&&&&&&&&#(/*,,,*//((((////(#&&&&&&&&&&&&&&&#((////////////(#&&&&&&#(*********//");
        $display(",***********,,,*,,*,,**************,,,*//******//(#&&&&&&&&&&&&&&&&&#(*,,*/(((#####(((((#&&&&&&&&&&&&&&&##///////////(#&&&&&&&&#(***///////");
        $display(",*************,,**,,,************,,,,,/(##((((####&&&&&&&&&&&&&&&&&&&(/**/(((#((((#((//(#&&&&&&&&&&&&&&&&&#(((((((((##&&&&&&&&&&#/**///////");
        $display(",******************************,,,,,,,*(#&#&&&&&&&&&&&&&&&&&&&&&&&&&&#(**/((#(#(((#((//(#&&&&&&&&&&&&&&&&&&&&&&&#&#&&&&&&&&&&&&&#(**///////");
        $display(",*************,**************,****,,,,,/(#&&&&&&&&&&&&&&&&&&&&&&&&&&&&#(/*/((((#((((///(#&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&(/*///////");
        $display(",*************************************,*/#&&&&&&&&&&&&&&&&&&&&&&&&&&&&&##(////////////(#&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&#/**/////*");
        $display(",******////****///////////////////////***/#&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&####(((((((###&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&#(********");
        $display(".,*,****///////////////////////////////***/#&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&#(/*******");
        $display(".,,,,*****//////////////////////////*******(#&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&##(*******");
        $display(".,,,,,,***********/////////////////********/(#&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&(*******");
        $display("=========================================");
    end
    else begin
        $display("Erorr number: %d", error_num);
        
        $display(" #######  ######   ######    #####   ######   ");
        $display("  ##   #   ##  ##   ##  ##  ##   ##   ##  ##  ");
        $display("  ## #     ##  ##   ##  ##  ##   ##   ##  ##  ");
        $display("  ####     #####    #####   ##   ##   #####   ");
        $display("  ## #     ## ##    ## ##   ##   ##   ## ##   ");
        $display("  ##   #   ##  ##   ##  ##  ##   ##   ##  ##  ");
        $display(" #######  #### ##  #### ##   #####   #### ##  ");
    end
    $finish;
end

initial begin
    #(`TOTAL_CYCLE);
    $display("Error : Time Out");
    $finish;
end

endmodule